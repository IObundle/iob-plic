`define iob_plic_ADDR_W 16