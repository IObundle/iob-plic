//add primary io to system instance
