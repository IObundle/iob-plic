//START_SWREG_TABLE clint
wire [`N_CORES-1:0] externalInterrupt;
